module uP_ROM
  #(
    parameter DATA_MAX_WIDTH = 29,
    parameter ADDR_WIDTH = 8
  ) (
    input wire [ADDR_WIDTH-1:0] addr,
    output wire [DATA_MAX_WIDTH-1:0] r_data
  );

  reg [DATA_MAX_WIDTH-1:0] u_ROM [0:2**ADDR_WIDTH-1];

  assign r_data = u_ROM[addr];

  initial begin
    //FETCH
    u_ROM[0] = 29'b00000010000001000000010110100;
    u_ROM[1] = 29'b00000000000001000000010000000;
    u_ROM[2] = 29'b01100000000010100000010000000;
    u_ROM[3] = 29'b00000000000000010001011000000;
    u_ROM[4] = 29'b00000000000000101000010000000;
    u_ROM[5] = 29'b01100010000010000011111000000;
    u_ROM[6] = 29'b00000000000000000000000000000;
    u_ROM[7] = 29'b00000000000000000000000000000;
	 //MOV A,ACC
	 u_ROM[8]  = 29'b10000011101110000001111000000;
    u_ROM[9]  = 29'b00000000000000000000000000000;
    u_ROM[10] = 29'b00000000000000000000000000000;
    u_ROM[11] = 29'b00000000000000000000000000000;
    u_ROM[12] = 29'b00000000000000000000000000000;
    u_ROM[13] = 29'b00000000000000000000000000000;
    u_ROM[14] = 29'b00000000000000000000000000000;
    u_ROM[15] = 29'b00000000000000000000000000000;
	 //MOV ACC,A
	 u_ROM[16] = 29'b10000001111110000001111000000;
    u_ROM[17] = 29'b00000000000000000000000000000;
    u_ROM[18] = 29'b00000000000000000000000000000;
    u_ROM[19] = 29'b00000000000000000000000000000;
    u_ROM[20] = 29'b00000000000000000000000000000;
    u_ROM[21] = 29'b00000000000000000000000000000;
    u_ROM[22] = 29'b00000000000000000000000000000;
    u_ROM[23] = 29'b00000000000000000000000000000;
	 //MOV ACC,CTE
	 u_ROM[24] = 29'b00000000000001000000010000000;
    u_ROM[25] = 29'b01100000000010100000010000000;
    u_ROM[26] = 29'b00000000011110010001111000000;
    u_ROM[27] = 29'b00000000000000000000000000000;
    u_ROM[28] = 29'b00000000000000000000000000000;
    u_ROM[29] = 29'b00000000000000000000000000000;
    u_ROM[30] = 29'b00000000000000000000000000000;
    u_ROM[31] = 29'b00000000000000000000000000000;
	 //MOV ACC,[DPTR]
	 u_ROM[32] = 29'b00000001000001000000010000000;
    u_ROM[33] = 29'b00000000000000110000010000000;
    u_ROM[34] = 29'b00000000011110010001111000000;
    u_ROM[35] = 29'b00000000000000000000000000000;
    u_ROM[36] = 29'b00000000000000000000000000000;
    u_ROM[37] = 29'b00000000000000000000000000000;
    u_ROM[38] = 29'b00000000000000000000000000000;
    u_ROM[39] = 29'b00000000000000000000000000000;
	 //MOV DPTR,ACC
	 u_ROM[40] = 29'b10000011101010000001111000000;
    u_ROM[41] = 29'b00000000000000000000000000000;
    u_ROM[42] = 29'b00000000000000000000000000000;
    u_ROM[43] = 29'b00000000000000000000000000000;
    u_ROM[44] = 29'b00000000000000000000000000000;
    u_ROM[45] = 29'b00000000000000000000000000000;
    u_ROM[46] = 29'b00000000000000000000000000000;
    u_ROM[47] = 29'b00000000000000000000000000000;
	 //MOV [DPTR],ACC
	 u_ROM[48] = 29'b00000001000001000000010000000;
    u_ROM[49] = 29'b10000011100000100000010000000;
    u_ROM[50] = 29'b00000000000000000011111000000;
    u_ROM[51] = 29'b00000000000000000000000000000;
    u_ROM[52] = 29'b00000000000000000000000000000;
    u_ROM[53] = 29'b00000000000000000000000000000;
    u_ROM[54] = 29'b00000000000000000000000000000;
    u_ROM[55] = 29'b00000000000000000000000000000;
	 //INV ACC
	 u_ROM[56] = 29'b10010011111110000001111000000;
    u_ROM[57] = 29'b00000000000000000000000000000;
    u_ROM[58] = 29'b00000000000000000000000000000;
    u_ROM[59] = 29'b00000000000000000000000000000;
    u_ROM[60] = 29'b00000000000000000000000000000;
    u_ROM[61] = 29'b00000000000000000000000000000;
    u_ROM[62] = 29'b00000000000000000000000000000;
    u_ROM[63] = 29'b00000000000000000000000000000;
	 //AND ACC,A
	 u_ROM[64] = 29'b10100001111110000001111000000;
    u_ROM[65] = 29'b00000000000000000000000000000;
    u_ROM[66] = 29'b00000000000000000000000000000;
    u_ROM[67] = 29'b00000000000000000000000000000;
    u_ROM[68] = 29'b00000000000000000000000000000;
    u_ROM[69] = 29'b00000000000000000000000000000;
    u_ROM[70] = 29'b00000000000000000000000000000;
    u_ROM[71] = 29'b00000000000000000000000000000;
	 //ADD ACC,A
	 u_ROM[72] = 29'b11010001111110000001111000000;
    u_ROM[73] = 29'b00000000000000000000000000000;
    u_ROM[74] = 29'b00000000000000000000000000000;
    u_ROM[75] = 29'b00000000000000000000000000000;
    u_ROM[76] = 29'b00000000000000000000000000000;
    u_ROM[77] = 29'b00000000000000000000000000000;
    u_ROM[78] = 29'b00000000000000000000000000000;
    u_ROM[79] = 29'b00000000000000000000000000000;
	 //JMP DIR
	 u_ROM[80] = 29'b00000000000001000000010000000;
    u_ROM[81] = 29'b00000000000000110000010000000;
    u_ROM[82] = 29'b00000000000010010001111000000;
    u_ROM[83] = 29'b00000000000000000000000000000;
    u_ROM[84] = 29'b00000000000000000000000000000;
    u_ROM[85] = 29'b00000000000000000000000000000;
    u_ROM[86] = 29'b00000000000000000000000000000;
    u_ROM[87] = 29'b00000000000000000000000000000;
	//JZ DIR
	 u_ROM[88] = 29'b00000000000001000000010010010;
    u_ROM[89] = 29'b01100000000010000001111000000;
    u_ROM[90] = 29'b00000000000000110000010000000;
    u_ROM[91] = 29'b00000000000010010001111000000;
    u_ROM[92] = 29'b00000000000000000000000000000;
    u_ROM[93] = 29'b00000000000000000000000000000;
    u_ROM[94] = 29'b00000000000000000000000000000;
    u_ROM[95] = 29'b00000000000000000000000000000;
	//JN DIR
	 u_ROM[96]  = 29'b00000000000001000000010011010;
    u_ROM[97]  = 29'b01100000000010000001111000000;
    u_ROM[98]  = 29'b00000000000000110000010000000;
    u_ROM[99]  = 29'b00000000000010010001111000000;
    u_ROM[100] = 29'b00000000000000000000000000000;
    u_ROM[101] = 29'b00000000000000000000000000000;
    u_ROM[102] = 29'b00000000000000000000000000000;
    u_ROM[103] = 29'b00000000000000000000000000000;
	//JC DIR
	 u_ROM[96]  = 29'b00000000000001000000010100010;
    u_ROM[97]  = 29'b01100000000010000001111000000;
    u_ROM[98]  = 29'b00000000000000110000010000000;
    u_ROM[99]  = 29'b00000000000010010001111000000;
    u_ROM[100] = 29'b00000000000000000000000000000;
    u_ROM[101] = 29'b00000000000000000000000000000;
    u_ROM[102] = 29'b00000000000000000000000000000;
    u_ROM[103] = 29'b00000000000000000000000000000;
	//SLL ACC
	 u_ROM[160] = 29'b10001011111110000001111000000;
    u_ROM[161] = 29'b00000000000000000000000000000;
    u_ROM[162] = 29'b00000000000000000000000000000;
    u_ROM[163] = 29'b00000000000000000000000000000;
    u_ROM[164] = 29'b00000000000000000000000000000;
    u_ROM[165] = 29'b00000000000000000000000000000;
    u_ROM[166] = 29'b00000000000000000000000000000;
    u_ROM[167] = 29'b00000000000000000000000000000;
	 //HALT
	 u_ROM[248] = 29'b00000000000000000000001000000;
    u_ROM[249] = 29'b00000000000000000000000000000;
    u_ROM[250] = 29'b00000000000000000000000000000;
    u_ROM[251] = 29'b00000000000000000000000000000;
    u_ROM[252] = 29'b00000000000000000000000000000;
    u_ROM[253] = 29'b00000000000000000000000000000;
    u_ROM[254] = 29'b00000000000000000000000000000;
    u_ROM[255] = 29'b00000000000000000000000000000;	 
  end

endmodule